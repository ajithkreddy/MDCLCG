module gpt(g, p, t, a, b);
output [63:0] g, p, t;
input [63:0] a,b;

and a0(g[0], a[0], b[0]);
or o0(p[0], a[0], b[0]);
xor x0(t[0], a[0], b[0]);

and a1(g[1], a[1], b[1]);
or o1(p[1], a[1], b[1]);
xor x1(t[1], a[1], b[1]);

and a2(g[2], a[2], b[2]);
or o2(p[2], a[2], b[2]);
xor x2(t[2], a[2], b[2]);

and a3(g[3], a[3], b[3]);
or o3(p[3], a[3], b[3]);
xor x3(t[3], a[3], b[3]);

and a4(g[4], a[4], b[4]);
or o4(p[4], a[4], b[4]);
xor x4(t[4], a[4], b[4]);

and a5(g[5], a[5], b[5]);
or o5(p[5], a[5], b[5]);
xor x5(t[5], a[5], b[5]);

and a6(g[6], a[6], b[6]);
or o6(p[6], a[6], b[6]);
xor x6(t[6], a[6], b[6]);

and a7(g[7], a[7], b[7]);
or o7(p[7], a[7], b[7]);
xor x7(t[7], a[7], b[7]);

and a8(g[8], a[8], b[8]);
or o8(p[8], a[8], b[8]);
xor x8(t[8], a[8], b[8]);

and a9(g[9], a[9], b[9]);
or o9(p[9], a[9], b[9]);
xor x9(t[9], a[9], b[9]);

and a10(g[10], a[10], b[10]);
or o10(p[10], a[10], b[10]);
xor x10(t[10], a[10], b[10]);

and a11(g[11], a[11], b[11]);
or o11(p[11], a[11], b[11]);
xor x11(t[11], a[11], b[11]);

and a12(g[12], a[12], b[12]);
or o12(p[12], a[12], b[12]);
xor x12(t[12], a[12], b[12]);

and a13(g[13], a[13], b[13]);
or o13(p[13], a[13], b[13]);
xor x13(t[13], a[13], b[13]);

and a14(g[14], a[14], b[14]);
or o14(p[14], a[14], b[14]);
xor x14(t[14], a[14], b[14]);

and a15(g[15], a[15], b[15]);
or o15(p[15], a[15], b[15]);
xor x15(t[15], a[15], b[15]);

and a16(g[16], a[16], b[16]);
or o16(p[16], a[16], b[16]);
xor x16(t[16], a[16], b[16]);

and a17(g[17], a[17], b[17]);
or o17(p[17], a[17], b[17]);
xor x17(t[17], a[17], b[17]);

and a18(g[18], a[18], b[18]);
or o18(p[18], a[18], b[18]);
xor x18(t[18], a[18], b[18]);

and a19(g[19], a[19], b[19]);
or o19(p[19], a[19], b[19]);
xor x19(t[19], a[19], b[19]);

and a20(g[20], a[20], b[20]);
or o20(p[20], a[20], b[20]);
xor x20(t[20], a[20], b[20]);

and a21(g[21], a[21], b[21]);
or o21(p[21], a[21], b[21]);
xor x21(t[21], a[21], b[21]);

and a22(g[22], a[22], b[22]);
or o22(p[22], a[22], b[22]);
xor x22(t[22], a[22], b[22]);

and a23(g[23], a[23], b[23]);
or o23(p[23], a[23], b[23]);
xor x23(t[23], a[23], b[23]);

and a24(g[24], a[24], b[24]);
or o24(p[24], a[24], b[24]);
xor x24(t[24], a[24], b[24]);

and a25(g[25], a[25], b[25]);
or o25(p[25], a[25], b[25]);
xor x25(t[25], a[25], b[25]);

and a26(g[26], a[26], b[26]);
or o26(p[26], a[26], b[26]);
xor x26(t[26], a[26], b[26]);

and a27(g[27], a[27], b[27]);
or o27(p[27], a[27], b[27]);
xor x27(t[27], a[27], b[27]);

and a28(g[28], a[28], b[28]);
or o28(p[28], a[28], b[28]);
xor x28(t[28], a[28], b[28]);

and a29(g[29], a[29], b[29]);
or o29(p[29], a[29], b[29]);
xor x29(t[29], a[29], b[29]);

and a30(g[30], a[30], b[30]);
or o30(p[30], a[30], b[30]);
xor x30(t[30], a[30], b[30]);

and a31(g[31], a[31], b[31]);
or o31(p[31], a[31], b[31]);
xor x31(t[31], a[31], b[31]);

and a32(g[32], a[32], b[32]);
or o32(p[32], a[32], b[32]);
xor x32(t[32], a[32], b[32]);

and a33(g[33], a[33], b[33]);
or o33(p[33], a[33], b[33]);
xor x33(t[33], a[33], b[33]);

and a34(g[34], a[34], b[34]);
or o34(p[34], a[34], b[34]);
xor x34(t[34], a[34], b[34]);

and a35(g[35], a[35], b[35]);
or o35(p[35], a[35], b[35]);
xor x35(t[35], a[35], b[35]);

and a36(g[36], a[36], b[36]);
or o36(p[36], a[36], b[36]);
xor x36(t[36], a[36], b[36]);

and a37(g[37], a[37], b[37]);
or o37(p[37], a[37], b[37]);
xor x37(t[37], a[37], b[37]);

and a38(g[38], a[38], b[38]);
or o38(p[38], a[38], b[38]);
xor x38(t[38], a[38], b[38]);

and a39(g[39], a[39], b[39]);
or o39(p[39], a[39], b[39]);
xor x39(t[39], a[39], b[39]);

and a40(g[40], a[40], b[40]);
or o40(p[40], a[40], b[40]);
xor x40(t[40], a[40], b[40]);

and a41(g[41], a[41], b[41]);
or o41(p[41], a[41], b[41]);
xor x41(t[41], a[41], b[41]);

and a42(g[42], a[42], b[42]);
or o42(p[42], a[42], b[42]);
xor x42(t[42], a[42], b[42]);

and a43(g[43], a[43], b[43]);
or o43(p[43], a[43], b[43]);
xor x43(t[43], a[43], b[43]);

and a44(g[44], a[44], b[44]);
or o44(p[44], a[44], b[44]);
xor x44(t[44], a[44], b[44]);

and a45(g[45], a[45], b[45]);
or o45(p[45], a[45], b[45]);
xor x45(t[45], a[45], b[45]);

and a46(g[46], a[46], b[46]);
or o46(p[46], a[46], b[46]);
xor x46(t[46], a[46], b[46]);

and a47(g[47], a[47], b[47]);
or o47(p[47], a[47], b[47]);
xor x47(t[47], a[47], b[47]);

and a48(g[48], a[48], b[48]);
or o48(p[48], a[48], b[48]);
xor x48(t[48], a[48], b[48]);

and a49(g[49], a[49], b[49]);
or o49(p[49], a[49], b[49]);
xor x49(t[49], a[49], b[49]);

and a50(g[50], a[50], b[50]);
or o50(p[50], a[50], b[50]);
xor x50(t[50], a[50], b[50]);

and a51(g[51], a[51], b[51]);
or o51(p[51], a[51], b[51]);
xor x51(t[51], a[51], b[51]);

and a52(g[52], a[52], b[52]);
or o52(p[52], a[52], b[52]);
xor x52(t[52], a[52], b[52]);

and a53(g[53], a[53], b[53]);
or o53(p[53], a[53], b[53]);
xor x53(t[53], a[53], b[53]);

and a54(g[54], a[54], b[54]);
or o54(p[54], a[54], b[54]);
xor x54(t[54], a[54], b[54]);

and a55(g[55], a[55], b[55]);
or o55(p[55], a[55], b[55]);
xor x55(t[55], a[55], b[55]);

and a56(g[56], a[56], b[56]);
or o56(p[56], a[56], b[56]);
xor x56(t[56], a[56], b[56]);

and a57(g[57], a[57], b[57]);
or o57(p[57], a[57], b[57]);
xor x57(t[57], a[57], b[57]);

and a58(g[58], a[58], b[58]);
or o58(p[58], a[58], b[58]);
xor x58(t[58], a[58], b[58]);

and a59(g[59], a[59], b[59]);
or o59(p[59], a[59], b[59]);
xor x59(t[59], a[59], b[59]);

and a60(g[60], a[60], b[60]);
or o60(p[60], a[60], b[60]);
xor x60(t[60], a[60], b[60]);

and a61(g[61], a[61], b[61]);
or o61(p[61], a[61], b[61]);
xor x61(t[61], a[61], b[61]);

and a62(g[62], a[62], b[62]);
or o62(p[62], a[62], b[62]);
xor x62(t[62], a[62], b[62]);

and a63(g[63], a[63], b[63]);
or o63(p[63], a[63], b[63]);
xor x63(t[63], a[63], b[63]);

endmodule
