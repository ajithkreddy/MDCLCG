module krgen(k, r, g, p);
output [63:0] k, r;
input [63:0] g, p;
wire w;

//k[0], r[0] to k[2], r[2]
assign k[0] = g[0];
assign r[0] = p[0];

or o0(k[1], g[1], g[0]);
and a0(r[1], p[1], p[0]);

and a1(w, p[1], g[0]);
or o1(k[2], g[2], g[1], w);
and a2(r[2], p[2], p[1], p[0]);


//k[3], r[3] to k[64], r[64]
kiri kr0(k[3], r[3], g[3:0], p[3:0]);
kiri kr1(k[4], r[4], g[4:1], p[4:1]);
kiri kr2(k[5], r[5], g[5:2], p[5:2]);
kiri kr3(k[6], r[6], g[6:3], p[6:3]);
kiri kr4(k[7], r[7], g[7:4], p[7:4]);

kiri kr5(k[8], r[8], g[8:5], p[8:5]);
kiri kr6(k[9], r[9], g[9:6], p[9:6]);
kiri kr7(k[10], r[10], g[10:7], p[10:7]);
kiri kr8(k[11], r[11], g[11:8], p[11:8]);
kiri kr9(k[12], r[12], g[12:9], p[12:9]);
kiri kr10(k[13], r[13], g[13:10], p[13:10]);
kiri kr11(k[14], r[14], g[14:11], p[14:11]);
kiri kr12(k[15], r[15], g[15:12], p[15:12]);

kiri kr13(k[16], r[16], g[16:13], p[16:13]);
kiri kr14(k[17], r[17], g[17:14], p[17:14]);
kiri kr15(k[18], r[18], g[18:15], p[18:15]);
kiri kr16(k[19], r[19], g[19:16], p[19:16]);
kiri kr17(k[20], r[20], g[20:17], p[20:17]);
kiri kr18(k[21], r[21], g[21:18], p[21:18]);
kiri kr19(k[22], r[22], g[22:19], p[22:19]);
kiri kr20(k[23], r[23], g[23:20], p[23:20]);

kiri kr21(k[24], r[24], g[24:21], p[24:21]);
kiri kr22(k[25], r[25], g[25:22], p[25:22]);
kiri kr23(k[26], r[26], g[26:23], p[26:23]);
kiri kr24(k[27], r[27], g[27:24], p[27:24]);
kiri kr25(k[28], r[28], g[28:25], p[28:25]);
kiri kr26(k[29], r[29], g[29:26], p[29:26]);
kiri kr27(k[30], r[30], g[30:27], p[30:27]);
kiri kr28(k[31], r[31], g[31:28], p[31:28]);

kiri kr29(k[32], r[32], g[32:29], p[32:29]);
kiri kr30(k[33], r[33], g[33:30], p[33:30]);
kiri kr31(k[34], r[34], g[34:31], p[34:31]);
kiri kr32(k[35], r[35], g[35:32], p[35:32]);
kiri kr33(k[36], r[36], g[36:33], p[36:33]);
kiri kr34(k[37], r[37], g[37:34], p[37:34]);
kiri kr35(k[38], r[38], g[38:35], p[38:35]);
kiri kr36(k[39], r[39], g[39:36], p[39:36]);

kiri kr37(k[40], r[40], g[40:37], p[40:37]);
kiri kr38(k[41], r[41], g[41:38], p[41:38]);
kiri kr39(k[42], r[42], g[42:39], p[42:39]);
kiri kr40(k[43], r[43], g[43:40], p[43:40]);
kiri kr41(k[44], r[44], g[44:41], p[44:41]);
kiri kr42(k[45], r[45], g[45:42], p[45:42]);
kiri kr43(k[46], r[46], g[46:43], p[46:43]);
kiri kr44(k[47], r[47], g[47:44], p[47:44]);

kiri kr45(k[48], r[48], g[48:45], p[48:45]);
kiri kr46(k[49], r[49], g[49:46], p[49:46]);
kiri kr47(k[50], r[50], g[50:47], p[50:47]);
kiri kr48(k[51], r[51], g[51:48], p[51:48]);
kiri kr49(k[52], r[52], g[52:49], p[52:49]);
kiri kr50(k[53], r[53], g[53:50], p[53:50]);
kiri kr51(k[54], r[54], g[54:51], p[54:51]);
kiri kr52(k[55], r[55], g[55:52], p[55:52]);

kiri kr53(k[56], r[56], g[56:53], p[56:53]);
kiri kr54(k[57], r[57], g[57:54], p[57:54]);
kiri kr55(k[58], r[58], g[58:55], p[58:55]);
kiri kr56(k[59], r[59], g[59:56], p[59:56]);
kiri kr57(k[60], r[60], g[60:57], p[60:57]);
kiri kr58(k[61], r[61], g[61:58], p[61:58]);
kiri kr59(k[62], r[62], g[62:59], p[62:59]);
kiri kr60(k[63], r[63], g[63:60], p[63:60]);

endmodule
