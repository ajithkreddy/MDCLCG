module Sgen(S, t, C);
output [63:0] S;
input [63:0] t;
input [63:0] C;

xor x0(S[0], t[0], C[0]);
xor x1(S[1], t[1], C[1]);
xor x2(S[2], t[2], C[2]);
xor x3(S[3], t[3], C[3]);
xor x4(S[4], t[4], C[4]);
xor x5(S[5], t[5], C[5]);
xor x6(S[6], t[6], C[6]);
xor x7(S[7], t[7], C[7]);

xor x8(S[8], t[8], C[8]);
xor x9(S[9], t[9], C[9]);
xor x10(S[10], t[10], C[10]);
xor x11(S[11], t[11], C[11]);
xor x12(S[12], t[12], C[12]);
xor x13(S[13], t[13], C[13]);
xor x14(S[14], t[14], C[14]);
xor x15(S[15], t[15], C[15]);

xor x16(S[16], t[16], C[16]);
xor x17(S[17], t[17], C[17]);
xor x18(S[18], t[18], C[18]);
xor x19(S[19], t[19], C[19]);
xor x20(S[20], t[20], C[20]);
xor x21(S[21], t[21], C[21]);
xor x22(S[22], t[22], C[22]);
xor x23(S[23], t[23], C[23]);

xor x24(S[24], t[24], C[24]);
xor x25(S[25], t[25], C[25]);
xor x26(S[26], t[26], C[26]);
xor x27(S[27], t[27], C[27]);
xor x28(S[28], t[28], C[28]);
xor x29(S[29], t[29], C[29]);
xor x30(S[30], t[30], C[30]);
xor x31(S[31], t[31], C[31]);

xor x32(S[32], t[32], C[32]);
xor x33(S[33], t[33], C[33]);
xor x34(S[34], t[34], C[34]);
xor x35(S[35], t[35], C[35]);
xor x36(S[36], t[36], C[36]);
xor x37(S[37], t[37], C[37]);
xor x38(S[38], t[38], C[38]);
xor x39(S[39], t[39], C[39]);

xor x40(S[40], t[40], C[40]);
xor x41(S[41], t[41], C[41]);
xor x42(S[42], t[42], C[42]);
xor x43(S[43], t[43], C[43]);
xor x44(S[44], t[44], C[44]);
xor x45(S[45], t[45], C[45]);
xor x46(S[46], t[46], C[46]);
xor x47(S[47], t[47], C[47]);

xor x48(S[48], t[48], C[48]);
xor x49(S[49], t[49], C[49]);
xor x50(S[50], t[50], C[50]);
xor x51(S[51], t[51], C[51]);
xor x52(S[52], t[52], C[52]);
xor x53(S[53], t[53], C[53]);
xor x54(S[54], t[54], C[54]);
xor x55(S[55], t[55], C[55]);

xor x56(S[56], t[56], C[56]);
xor x57(S[57], t[57], C[57]);
xor x58(S[58], t[58], C[58]);
xor x59(S[59], t[59], C[59]);
xor x60(S[60], t[60], C[60]);
xor x61(S[61], t[61], C[61]);
xor x62(S[62], t[62], C[62]);
xor x63(S[63], t[63], C[63]);

endmodule
